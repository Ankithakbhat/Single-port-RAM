 `include "ram_trx.sv"
 `include "ram_gen.sv"
 `include "ram_drv.sv"
 `include "ram_moni.sv"
 `include "ram_ref_model.sv"
 `include "ram_sb.sv"
 `include "ram_env.sv"
 `include "ram_test.sv"
`include "interface.sv"
